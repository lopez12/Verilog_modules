`timescale 1ns/100ps
module AsyncSimpleLogic_top
(    
    output  [6:0]   seg,
    output  dp,

    output  [3:0]   an,

    output  [7:0]   Led,

    input   [7:0]   sw,

    input   [3:0]   btn
);


//
//----------------------------------------------------------------------------------
//
// Start of test achitecture
//
//
//----------------------------------------------------------------------------------
	// --------------------------------------------------------------------------
	//                        Continuous Assignments
	// --------------------------------------------------------------------------

	assign	Led[0]		    =		btn[0];
	assign	Led[1]		    =		~btn[1];
	assign	Led[2]		    =		btn[0] & btn[1];
	assign	Led[3]		    =		btn[0] | btn[1];
	assign	Led[4]		    =		~(btn[0] & btn[1]);
	assign	Led[5]		    =		~(btn[0] | btn[1]);
	assign	Led[6]		    =		btn[0] ^ btn[1];
	assign	Led[7]		    =		~(btn[0] ^ btn[1]);

	assign	seg[6:0]		=		sw[6:0];
	assign	dp				=		~sw[7];
	assign	an[0]			=		btn[2]|btn[3];
	assign	an[1]			=		btn[2]|~btn[3];
	assign	an[2]			=		~btn[2]|btn[3];
	assign	an[3]			=		~(btn[2]&btn[3]);
	
//----------------------------------------------------------------------------------------------------------------------------------------------------------------------
//
// Start of circuit description
//
endmodule
// --------------------------------------------------------------------------
//                    End Of File              
// --------------------------------------------------------------------------
